* Title: Passive RL LPF

* Netlist
Vin 1 0 dc 0 ac 1
L1 1 2 159m
R1 2 0 10k
.end
