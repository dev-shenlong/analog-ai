* Title: Parallel R

* Netlist:
Vin 1 0 dc 1
R1 1 0 1k
R2 1 0 2k
R3 1 0 3k
.end
